`ifndef __DEC_CONFIGS_SV
`define __DEC_CONFIGS_SV


//  Package: ncu_configs
//
package configs;

  //  Group: Parameters
  localparam unsigned LiftingFactor = 81;
  localparam unsigned DWIDTH = 5;

endpackage : configs

`endif
